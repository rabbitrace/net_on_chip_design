
module hex (
	probe);	

	input	[30:0]	probe;
endmodule
